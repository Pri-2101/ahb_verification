
package env_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    import apb_slave_agent_pkg::*;
    import apb_master_agent_pkg::*;

    `include "env_config.svh"
    `include "env.svh"
    `include "apb_master_single_trans_sequence.svh"
    `include "apb_master_INCR_sequence.svh"
    `include "apb_slave_single_trans_sequence.svh"
    `include "apb_master_complete_sequence.svh"

endpackage : env_pkg
