package apb_slave_agent_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"
`include "param_enums.svh"

//import register_layering_pkg::*;
//`include "apb_monitor_assertions.svh"
`include "apb_slave_seq_item.svh"
`include "apb_slave_agent_config.svh"
`include "apb_slave_driver.svh"
`include "apb_slave_monitor.svh"
`include "apb_slave_sequencer.svh"
//`include "apb_listener.svh"
`include "apb_slave_agent.sv"


// Utility Sequences
//`include "apb_slave_sequence.svh"

endpackage: apb_slave_agent_pkg
